`timescale 1ns / 1ps

module top
(
    input                                   i_reset,
    input                                   i_clock,
    input                                   i_serial_start,
    output                                  o_serial
);  
    
    /* System */
    wire            clock;
    wire            locked;
    
    /* Serial */
    localparam  SERIAL_DATA_SIZE    =   8;
    
    /* ADC */
    localparam  ADC_DATA_SIZE       =   16;
    wire                                    adc_clock;
    
    /* ###################################### */
    clk_wiz_0
    u_clk_wiz_0
    (
        .clk_in1                (i_clock),
        .reset                  (i_reset),
        .clk_out1               (clock),
        .clk_out2               (adc_clock),
        .locked                 (locked)
    );
    /* ###################################### */
    serial #
    (
        .SERIAL_DATA_SIZE       (SERIAL_DATA_SIZE)
    )
    u_serial
    (
        .i_clock                (clock),
        .i_reset                (~locked),
        .i_start                (i_serial_start),
        .o_serial               (o_serial)
    );
    /* ###################################### */
    /*
    ZmodADC1410_Controller_0
    u_ZmodADC1410_Controller_0
    (
        .SysClk     (clock),
        .ADC_InClk  (adc_clock),
        .sRst_n     (~locked),
        .sCh1Out    (tx_data)
    );
    */
    /* ###################################### */

endmodule


/*
    SysClk :        IN STD_LOGIC;                          100mhz input clock
    ADC_InClk :     IN STD_LOGIC;                       400mhz input clock
    sRst_n :        IN STD_LOGIC;                          synchronous reset negative polarity
    sInitDone_n :       OUT STD_LOGIC;                    active low flag, inidicate zmod initialization complete
    FIFO_EMPTY_CHA :    OUT STD_LOGIC;                 
    FIFO_EMPTY_CHB :    OUT STD_LOGIC;
    sCh1Out :           OUT STD_LOGIC_VECTOR(15 DOWNTO 0);    output data ch1 synchronoues with sysclk
    sTestMode :     IN STD_LOGIC;                       
    adcClkIn_p :        OUT STD_LOGIC;                     adc positive differential clock input
    adcClkIn_n :        OUT STD_LOGIC;                     adc negative differential clock input
    adcSync :           OUT STD_LOGIC;                        synchronitazino signal
    DcoClk :        IN STD_LOGIC;                          data strobe generated by the ADC used to captura dADC_Data
    dADC_Data :     IN STD_LOGIC_VECTOR(13 DOWNTO 0);   ddr parallel data bus exportes by ADC containgin ch1 and ch2 multiplexed samples
    sADC_SDIO :             INOUT STD_LOGIC;                    spi sdio signal
    sADC_CS :           OUT STD_LOGIC;                        spi cs signal
    sADC_Sclk :         OUT STD_LOGIC;                      spi output clock
    sCh1CouplingH :     OUT STD_LOGIC;                  Channel1 AC DC coupling relay driver control input.
    sCh1CouplingL :     OUT STD_LOGIC;                  Channel1 AC DC coupling select relay driver control input
    sCh1GainH :         OUT STD_LOGIC;                      Channel1 gain select relay driver control input.
    sCh1GainL :         OUT STD_LOGIC;                      Channel1 gain select relay driver control input.
    sRelayComH :        OUT STD_LOGIC;                     Common relay terminal driver control input.
    sRelayComL :        OUT STD_LOGIC                      Common relay terminal driver control input.
    
    sExtCh1LgMultCoef :     IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    sExtCh1LgAddCoef :      IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    sExtCh1HgMultCoef :     IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    sExtCh1HgAddCoef :      IN STD_LOGIC_VECTOR(17 DOWNTO 0);
*/